Ripple problem
Vin 3 1 sin(0,15,50,0,0)
D1 1 2 diode1
D2 3 2 diode2
D3 0 3 diode3
D4 0 1 diode4
.model diode1 D
.model diode2 D
.model diode3 D
.model diode4 D
C1 2 0 44.4u
R1 2 0 500 1500
.control
tran 0.0000001 40m
set color0 = white
set color1 = black
set color1 = blue
plot tran.v(2) 
.endc
.end
